module bus(
    
);


    
endmodule