module master_mux(
    port_list
);
    
endmodule